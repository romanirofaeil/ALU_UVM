package alu_package;
    import uvm_pkg::*;
    `include "alu_sequence_item.sv"
    `include "alu_sequence_config.sv"
    `include "alu_sequence.sv"
    `include "alu_ADD_sequence.sv"
    `include "alu_SUB_sequence.sv"
    `include "alu_XOR_sequence.sv"
    `include "alu_AND_sequence.sv"
    `include "alu_OR_sequence.sv"
    `include "alu_XNOR_sequence.sv"
    `include "alu_NAND_sequence.sv"
    `include "alu_A_MINUS_1_sequence.sv"
    `include "alu_B_PLUS_2_sequence.sv"
    `include "alu_ERROR_sequence.sv"
    `include "alu_sequencer.sv"
    `include "alu_agent_config.sv"
    `include "alu_driver.sv"
    `include "alu_monitor.sv"
    `include "alu_agent.sv"
    `include "alu_scoreboard.sv"
    `include "alu_functional_coverage.sv"
    `include "alu_environment.sv"
    `include "alu_test.sv"
    `include "alu_ADD_test.sv"
    `include "alu_SUB_test.sv"
    `include "alu_XOR_test.sv"
    `include "alu_AND_test.sv"
    `include "alu_OR_test.sv"
    `include "alu_XNOR_test.sv"
    `include "alu_NAND_test.sv"
    `include "alu_A_MINUS_1_test.sv"
    `include "alu_B_PLUS_2_test.sv"
    `include "alu_ERORR_test.sv"
endpackage
